module ControlUnitOutput(
	input [5:0] OPCode, 
	input [2:0] CurrentState, 
	output reg [54:0] ControlSignals);
	
	always@(*)
	begin
		case(CurrentState)
			3'b000: //First cycle control signals
				begin
					ControlSignals[0] = 1'b1; //PCRead;
					ControlSignals[1] = 1'b0; //IRWrite;
					ControlSignals[3:2] = 2'bxx; //MUXULAInp1Select;
					ControlSignals[5:4] = 2'bxx; //MUXULAInp2Select;
					ControlSignals[7:6] = 2'bxx; //MUXULAInp3Select;
					ControlSignals[8] = 1'bx; //MUXPCInpSelect;
					ControlSignals[10:9] = 2'b01; //AddressMUXSelect;
					ControlSignals[11] = 1'b0; //AddressRead;
					ControlSignals[12] = 1'b0; //MemDataRead;
					ControlSignals[13] = 1'b0; //PCWrite;
					ControlSignals[14] = 1'b0; //IRRead;
					ControlSignals[15] = 1'b0; //AccRead;
					ControlSignals[16] = 1'b0; //AccWrite;
					ControlSignals[17] = 1'b0; //SPRead;
					ControlSignals[18] = 1'b0; //SPWrite;
					ControlSignals[19] = 1'b0; //XRead;
					ControlSignals[20] = 1'b0; //XWrite;
					ControlSignals[21] = 1'b0; //YRead;
					ControlSignals[22] = 1'b0; //YWrite;
					ControlSignals[25:23] = 3'bxxx; //ULAControl;
					ControlSignals[27:26] = 2'bxx; //MemWriteSelect;
					ControlSignals[29:28] = 2'bxx; //MemWriteSelect2;
					ControlSignals[30] = 1'b0; //MemDataWrite;
					ControlSignals[31] = 1'b0; //ProcessorStatusRead;
					ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
					ControlSignals[33] = 1'b0; //ALURead;
					ControlSignals[34] = 1'bx; //MUXPCInp2Select;
					ControlSignals[38:35] = 4'b0000; //BranchSignals;
					ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
					ControlSignals[44:42] = 3'b000; //SRClearsSignals;
					ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b1; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
				end
			3'b001: //Second cycle control signals
				begin
					ControlSignals[0] = 1'b0; //PCRead;
					ControlSignals[1] = 1'b1; //IRWrite;
					ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
					ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
					ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
					ControlSignals[8] = 1'b0; //MUXPCInpSelect;
					ControlSignals[10:9] = 2'b01; //AddressMUXSelect;
					ControlSignals[11] = 1'b0; //AddressRead;
					ControlSignals[12] = 1'b1; //MemDataRead;
					ControlSignals[13] = 1'b1; //PCWrite;
					ControlSignals[14] = 1'b0; //IRRead;
					ControlSignals[15] = 1'b0; //AccRead;
					ControlSignals[16] = 1'b0; //AccWrite;
					ControlSignals[17] = 1'b0; //SPRead;
					ControlSignals[18] = 1'b0; //SPWrite;
					ControlSignals[19] = 1'b0; //XRead;
					ControlSignals[20] = 1'b0; //XWrite;
					ControlSignals[21] = 1'b0; //YRead;
					ControlSignals[22] = 1'b0; //YWrite;
					ControlSignals[25:23] = 3'b000; //ULAControl;
					ControlSignals[27:26] = 2'bxx; //MemWriteSelect;
					ControlSignals[29:28] = 2'bxx; //MemWriteSelect2;
					ControlSignals[30] = 1'b0; //MemDataWrite;
					ControlSignals[31] = 1'b0; //ProcessorStatusRead;
					ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
					ControlSignals[33] = 1'b1; //ALURead;
					ControlSignals[34] = 1'b0; //MUXPCInp2Select;
					ControlSignals[38:35] = 4'b0000; //BranchSignals;
					ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
					ControlSignals[44:42] = 3'b000; //SRClearsSignals;
					ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
				end
			3'b010: //Third cycle control signals
				begin
					ControlSignals[0] = 1'b0; //PCRead;
					ControlSignals[1] = 1'b0; //IRWrite;
					ControlSignals[3:2] = 2'bxx; //MUXULAInp1Select;
					ControlSignals[5:4] = 2'bxx; //MUXULAInp2Select;
					ControlSignals[7:6] = 2'bxx; //MUXULAInp3Select;
					ControlSignals[8] = 1'b0; //MUXPCInpSelect;
					ControlSignals[10:9] = 2'b10; //AddressMUXSelect;
					ControlSignals[11] = 1'b0; //AddressRead;
					ControlSignals[12] = 1'b0; //MemDataRead;
					ControlSignals[13] = 1'b0; //PCWrite;
					ControlSignals[14] = 1'b0; //IRRead;
					ControlSignals[15] = 1'b0; //AccRead;
					ControlSignals[16] = 1'b0; //AccWrite;
					ControlSignals[17] = 1'b0; //SPRead;
					ControlSignals[18] = 1'b0; //SPWrite;
					ControlSignals[19] = 1'b0; //XRead;
					ControlSignals[20] = 1'b0; //XWrite;
					ControlSignals[21] = 1'b0; //YRead;
					ControlSignals[22] = 1'b0; //YWrite;
					ControlSignals[25:23] = 3'bxxx; //ULAControl;
					ControlSignals[27:26] = 2'bxx; //MemWriteSelect;
					ControlSignals[29:28] = 2'bxx; //MemWriteSelect2;
					ControlSignals[30] = 1'b0; //MemDataWrite;
					ControlSignals[31] = 1'b0; //ProcessorStatusRead;
					ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
					ControlSignals[33] = 1'b0; //ALURead;
					ControlSignals[34] = 1'b0; //MUXPCInp2Select;
					ControlSignals[38:35] = 4'b0000; //BranchSignals;
					ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
					ControlSignals[44:42] = 3'b000; //SRClearsSignals;
					ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
				end
			3'b011: //Fourth cycle control signals
				case(OPCode)
					6'b000000: //CPY
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b1; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b000001: //CPI
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b1; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b000010: //CMP
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b1; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b000011: //ASL
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b010; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b000100: //ANDI
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b001; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b000101: //AND
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b001; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b000110: //ADCI
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b000111: //ADC
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
						6'b001000: //TXAX
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b1; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b01; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b001001: //SBCI
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b001010: //SBC
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b001011: //ORAI
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b110; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b001100: //ORA
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b110; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b001101: //LSR
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b101; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b001110: //EORI
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b100; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b001111: //EOR
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b100; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b010000: //TAXX
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b1; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b10; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b010001: //STA
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b1; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b10; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b101; //ULAControl;
							ControlSignals[27:26] = 2'b10; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b1; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b010010: //LDYI
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b10; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b10; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b1; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b010011: //LDY
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b10; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b10; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b1; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b010100: //LDXI
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b10; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b10; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b1; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
							ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b010101: //LDX
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b10; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b10; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b1; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
							ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b010110: //LDAI
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b10; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b10; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b010111: //LDA
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b10; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b10; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011000: //TAXBR
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b10; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b1; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b10; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011001: //TXS
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b10; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b1; //SPWrite;
							ControlSignals[19] = 1'b1; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011010: //TSX
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b10; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b1; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b1; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011011: //PLP
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b10; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b1; //AddressRead;
							ControlSignals[12] = 1'b1; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b1; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011100: //PLA
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b101; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b1; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011101: //PHP
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b1; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b01; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011110: //PHA
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b1; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011111: //STY
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b1; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b10; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b101; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b1; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
						6'b100000: //PHPC
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b1; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b100001: //RTS
						begin 
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b101; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b1; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b100010: //JSR
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b1; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b100011: //JMP
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b1; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b1; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b101; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b100100: //BPL
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b1; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0001; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b100101: //BNE
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b1; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0010; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b100110: //BMI
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b1; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0100; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b100111: //BEQ
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b1; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b1000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
						6'b101000: //PLPC
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b101; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b1; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
							ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b110000: //TYA
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b1; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b110001: //TXA
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b1; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b110010: //TAY
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b1; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b1; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b110011: //TAX
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b1; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b1; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b110100: //INY
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b1; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b110101: //INX
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b1; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
					ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b110110: //DEY
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b10; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b1; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b110111: //DEX
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b1; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
						6'b111000: //SPC
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b1; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b1; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b10; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
							ControlSignals[54] = 1'b1; //savedPCReadSignal;
						end
					6'b111001: //SFF
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b1; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b1; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
						6'b111010: //CPF
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b1; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b1; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b111100: //INT
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b01; //OutputInputSignal;
							ControlSignals[41] = 1'b1; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b111011: //OUP
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b10; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b101001: //DIVI
					begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b1; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
					end
					6'b101010: //DIV
					begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b1; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
					end
					6'b101011: //MULI
					begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b11; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b1; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
					end
					6'b101100: //MUL
					begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b1; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
							
					end
					6'b101101: //CLV
					begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b001; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b101110: //CLN
					begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b010; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
					end
					6'b101111: //CLZ
					begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b100; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
					end
					6'b111110: //NOP
					begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
					end
					6'b111111: //BRK
					begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b1; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
					end
					default:
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
					ControlSignals[46] = 1'b0; //ALUExtra;
					ControlSignals[47] = 1'b0; //BRWriteSignal;
					ControlSignals[48] = 1'b0; //CountSignal;
					ControlSignals[49] = 1'b0; //CFFSignal;
					ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					endcase
			3'b100: //Fifth cycle control signals
				case(OPCode)
					6'b011011: //PLP
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b1; //AddressRead;
							ControlSignals[12] = 1'b1; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b1; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b1; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011100: //PLA
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b1; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b1; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b1; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011101: //PHP
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b1; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b10; //MemWriteSelect;
							ControlSignals[29:28] = 2'b01; //MemWriteSelect2;
							ControlSignals[30] = 1'b1; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b011110: //PHA
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b1; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b10; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b1; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
						6'b100000: //PHPC
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b11; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b1; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
							ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b101000: //PLPC
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b1; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b1; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b1; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
							ControlSignals[53] = 1'b1; //savedPCWriteSignal;
							ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b100001: //RTS
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b1; //MemDataRead;
							ControlSignals[13] = 1'b1; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b1; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b1; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b100010: //JSR
						begin
							ControlSignals[0] = 1'b1; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b01; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b10; //MemWriteSelect;
							ControlSignals[29:28] = 2'b10; //MemWriteSelect2;
							ControlSignals[30] = 1'b1; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
							ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b111100: //INT
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b1; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b01; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					6'b111111: //BRK
					begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b1; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
					end
					default:
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b01; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b1; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b011; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
				endcase
			3'b101: //Sixth cycle control signals
				case(OPCode)
					6'b100010: //JSR
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b11; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b01; //MUXULAInp3Select;
							ControlSignals[8] = 1'b1; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b1; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b101; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b1; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					default:
						begin
							ControlSignals[0] = 1'b0; //PCRead;
							ControlSignals[1] = 1'b0; //IRWrite;
							ControlSignals[3:2] = 2'b00; //MUXULAInp1Select;
							ControlSignals[5:4] = 2'b00; //MUXULAInp2Select;
							ControlSignals[7:6] = 2'b00; //MUXULAInp3Select;
							ControlSignals[8] = 1'b0; //MUXPCInpSelect;
							ControlSignals[10:9] = 2'b00; //AddressMUXSelect;
							ControlSignals[11] = 1'b0; //AddressRead;
							ControlSignals[12] = 1'b0; //MemDataRead;
							ControlSignals[13] = 1'b0; //PCWrite;
							ControlSignals[14] = 1'b0; //IRRead;
							ControlSignals[15] = 1'b0; //AccRead;
							ControlSignals[16] = 1'b0; //AccWrite;
							ControlSignals[17] = 1'b0; //SPRead;
							ControlSignals[18] = 1'b0; //SPWrite;
							ControlSignals[19] = 1'b0; //XRead;
							ControlSignals[20] = 1'b0; //XWrite;
							ControlSignals[21] = 1'b0; //YRead;
							ControlSignals[22] = 1'b0; //YWrite;
							ControlSignals[25:23] = 3'b000; //ULAControl;
							ControlSignals[27:26] = 2'b00; //MemWriteSelect;
							ControlSignals[29:28] = 2'b00; //MemWriteSelect2;
							ControlSignals[30] = 1'b0; //MemDataWrite;
							ControlSignals[31] = 1'b0; //ProcessorStatusRead;
							ControlSignals[32] = 1'b0; //ProcessorStatusWrite;
							ControlSignals[33] = 1'b0; //ALURead;
							ControlSignals[34] = 1'b0; //MUXPCInp2Select;
							ControlSignals[38:35] = 4'b0000; //BranchSignals;
							ControlSignals[40:39] = 2'b00; //OutputInputSignal;
							ControlSignals[41] = 1'b0; //WaitingInput;
							ControlSignals[44:42] = 3'b000; //SRClearsSignals;
							ControlSignals[45] = 1'b0; //BRKSignal;
							ControlSignals[46] = 1'b0; //ALUExtra;
							ControlSignals[47] = 1'b0; //BRWriteSignal;
							ControlSignals[48] = 1'b0; //CountSignal;
							ControlSignals[49] = 1'b0; //CFFSignal;
							ControlSignals[50] = 1'b0; //procFinishSignal;
					ControlSignals[52:51] = 2'b00; //AuxSignals;
					ControlSignals[53] = 1'b0; //savedPCWriteSignal;
					ControlSignals[54] = 1'b0; //savedPCReadSignal;
						end
					endcase
				default: ControlSignals = 46'd0;
		endcase
	end

endmodule
